LIBRARY ieee; 
USE ieee.std_logic_1164.all;

ENTITY latch2 IS 
	PORT (A : IN STD_LOGIC_VECTOR(7 DOWNTO 0); --8 BIT A INPUT
			RESET, CLOCK: IN STD_LOGIC; -- 1 BIT CLOCK AND RESET
			Q: OUT STD_LOGIC_VECTOR (7 DOWNTO 0));-- 8 BIT Q OUTPUT
END latch2; 
ARCHITECTURE BEHAVIOR OF latch2 IS
BEGIN 
	PROCESS (RESET, CLOCK)
	BEGIN
		IF RESET = '0' THEN Q <= "00000000"; 
		ELSIF CLOCK'EVENT AND CLOCK = '0'THEN Q<=A;
		END IF;
	END PROCESS;
END BEHAVIOR;