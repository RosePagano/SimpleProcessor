LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY ALUcore IS 
PORT( CLOCK: IN STD_LOGIC;
		A, B: IN UNSIGNED(7 DOWNTO 0);
		OP: IN UNSIGNED(15 DOWNTO 0);
		NEG: OUT STD_LOGIC;
		R1, R2: OUT UNSIGNED(3 DOWNTO 0));
END ALUcore; 
ARCHITECTURE CALCULATION OF ALUcore IS 
SIGNAL REG1, REG2, RESULT: UNSIGNED(7 DOWNTO 0):=(OTHERS => '0');
SIGNAL REG4: UNSIGNED(0 DOWNTO 7);
BEGIN
REG1 <=A;
REG2 <=B;
PROCESS(CLOCK, OP)
BEGIN
	IF(RISING_EDGE(CLOCK)) THEN 
		CASE OP IS 
			WHEN "0000000000000001" => --ADD 
			NEG <= '0';
			RESULT <= (REG1 + REG2);
			WHEN "0000000000000010" =>  --SUBTRACT
				IF(REG1 >= REG2) THEN 
					RESULT <= (REG1 - REG2); 
					NEG <= '0';
				ELSE 
					NEG <= '1'; 
					RESULT <= (REG2 - REG1);
				END IF;
			WHEN "0000000000000100" => RESULT <= NOT(REG1);--NOT
			WHEN "0000000000001000" => RESULT <= NOT(REG1 AND REG2); --NOT (A AND B)
			WHEN "0000000000010000" => RESULT <= NOT(REG1 OR REG2);--NOT (A OR B)
			WHEN "0000000000100000" => RESULT <= REG1 AND REG2;--A AND B
			WHEN "0000000001000000" => RESULT <= REG1 XOR REG2; --A XOR B
			WHEN "0000000010000000" => RESULT <= REG1 OR REG2;--A OR B
			WHEN "0000000100000000" => RESULT <= NOT(REG1 XOR REG2); --NOT(A XOR B)
			WHEN OTHERS => -- DO NOTHING
			RESULT <= "00000000";
		END CASE;
	END IF;
END PROCESS;
R1 <= RESULT(3 DOWNTO 0);
R2 <= RESULT(7 DOWNTO 4);
end calculation; 