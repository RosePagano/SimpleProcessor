LIBRARY ieee; 
USE ieee.std_logic_1164.all;

ENTITY ADD IS 
	PORT (OP1, OP2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0); --8 BIT A INPUT
			OPOUT: OUT STD_LOGIC_VECTOR (15 DOWNTO 0));-- 8 BIT Q OUTPUT
END ADD; 
ARCHITECTURE BEHAVIOR OF ADD IS
BEGIN 
	PROCESS (OP1, OP2)
	BEGIN
		OPOUT <= OP1(7 DOWNTO 0);
		OPOUT <= OP2(15 DOWNTO 8);
	END PROCESS;
END BEHAVIOR;