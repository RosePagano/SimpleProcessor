LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY decod4to16 IS 
	PORT (W : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			En : IN STD_LOGIC;
			Y : OUT STD_LOGIC_VECTOR(15 DOWNTO 0));
END decod4to16; 

ARCHITECTURE Behavior OF decod4to16 IS
BEGIN
	PROCESS (W,En)
BEGIN
	IF (En = '0') THEN
	Y <= "0000000000000000";
	ELSE
	CASE W is
		WHEN "0000" =>
		 Y <= "0000000000000001";
		WHEN "0001" =>
		 Y <= "0000000000000010";
		WHEN "0010" =>
		 Y <= "0000000000000100";
		WHEN "0011" =>
		 Y <= "0000000000001000";
		WHEN "0100" =>
		 Y <= "0000000000010000";
		WHEN "0101" =>
		 Y <= "0000000000100000";
		WHEN "0110" =>
		 Y <= "0000000001000000";
		WHEN "0111" =>
		 Y <= "0000000010000000";
		WHEN "1000" =>
		 Y <= "0000000100000000";
		WHEN "1001" =>
		 Y <= "0000001000000000";
		WHEN "1010" =>
		 Y <= "0000010000000000";
		WHEN "1011" =>
		 Y <= "0000100000000000";
		WHEN "1100" =>
		 Y <= "0001000000000000";
		WHEN "1101" =>
		 Y <= "0010000000000000";
		WHEN "1110" =>
		 Y <= "0100000000000000";
		WHEN "1111" =>
		 Y <= "1000000000000000";
	WHEN OTHERS => Y <= "0000000000000000";
	END CASE;
END IF;
END PROCESS;
END behavior;	